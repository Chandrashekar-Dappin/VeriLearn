//demo file

module demo;
endmodule
